`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    18:12:10 11/06/2012 
// Design Name: 
// Module Name:    FPGATop 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module FPGATop(
   input clk, 
   input [7:0] Qie1_Out,Qie2_Out,Qie3_Out,Qie4_Out,
               Qie5_Out,Qie6_Out,Qie7_Out,Qie8_Out,
               Qie9_Out,Qie10_Out,Qie11_Out,Qie12_Out,
   input       Qie1_CkOut,Qie2_CkOut,Qie3_CkOut,Qie4_CkOut,
               Qie5_CkOut,Qie6_CkOut,Qie7_CkOut,Qie8_CkOut,
               Qie9_CkOut,Qie10_CkOut,Qie11_CkOut,Qie12_CkOut,
   input       Qie1_DiscOut,Qie2_DiscOut,Qie3_DiscOut,Qie4_DiscOut,
               Qie5_DiscOut,Qie6_DiscOut,Qie7_DiscOut,Qie8_DiscOut,
               Qie9_DiscOut,Qie10_DiscOut,Qie11_DiscOut,Qie12_DiscOut
   );

endmodule
